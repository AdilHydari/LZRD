MFB_BANDPASS.CIR - OPAMP MULTIPLE FEEDBACK BAND-PASS FILTER
*

VS	1	0	AC	1	SIN(0VOFF  1VPEAK 10KHZ)
*
R1A	1	2	7.96K
R1B	2	0	162
R2	3	4	15.9K
C1	2	3	10000PF
C2	2	4	10000PF
*
XOP	0	3 4	OPAMP1
*
*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
* GBP = DCGAIN X POLE1 = 10MHz
EGAIN   3 0     1 2     100K
RP1     3       4       1000
CP1     4       0       1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER 5 0     4 0     1
ROUT    5       6       10
.ENDS
*
* ANALYSIS
.AC 	DEC 	200 3K 30K
*.TRAN	1US 1000US
*
* VIEW RESULTS
.PROBE
.END
